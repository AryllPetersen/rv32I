`include "rv32I.h"


module ControlUnit(
  input logic clock, resetn,
  input logic[31:0] ir,
  input irsel_t irsel,
  input pcsel_t pcsel,
  

);


endmodule